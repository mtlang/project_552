module Decoder_7_128(tag, block);

input [6:0] tag;

output [127:0] block;

assign block = (tag == 0) ? 128'h00000000000000000000000000000000 :
				(tag == 1) ? 128'h00000000000000000000000000000001 :
				(tag == 2) ? 128'h00000000000000000000000000000002 :
				(tag == 3) ? 128'h00000000000000000000000000000004 :
				(tag == 4) ? 128'h00000000000000000000000000000008 :
				(tag == 5) ? 128'h00000000000000000000000000000010 :
				(tag == 6) ? 128'h00000000000000000000000000000020 :
				(tag == 7) ? 128'h00000000000000000000000000000040 :
				(tag == 8) ? 128'h00000000000000000000000000000080 :
				(tag == 9) ? 128'h00000000000000000000000000000100 :
				(tag == 10) ? 128'h00000000000000000000000000000200 :
				(tag == 11) ? 128'h00000000000000000000000000000400 :
				(tag == 12) ? 128'h00000000000000000000000000000800 :
				(tag == 13) ? 128'h00000000000000000000000000001000 :
				(tag == 14) ? 128'h00000000000000000000000000002000 :
				(tag == 15) ? 128'h00000000000000000000000000004000 :
				(tag == 16) ? 128'h00000000000000000000000000008000 :
				(tag == 17) ? 128'h00000000000000000000000000010000 :
				(tag == 18) ? 128'h00000000000000000000000000020000 :
				(tag == 19) ? 128'h00000000000000000000000000040000 :
				(tag == 20) ? 128'h00000000000000000000000000080000 :
				(tag == 21) ? 128'h00000000000000000000000000100000 :
				(tag == 22) ? 128'h00000000000000000000000000200000 :
				(tag == 23) ? 128'h00000000000000000000000000400000 :
				(tag == 24) ? 128'h00000000000000000000000000800000 :
				(tag == 25) ? 128'h00000000000000000000000001000000 :
				(tag == 26) ? 128'h00000000000000000000000002000000 :
				(tag == 27) ? 128'h00000000000000000000000004000000 :
				(tag == 28) ? 128'h00000000000000000000000008000000 :
				(tag == 29) ? 128'h00000000000000000000000010000000 :
				(tag == 30) ? 128'h00000000000000000000000020000000 :
				(tag == 31) ? 128'h00000000000000000000000040000000 :
				(tag == 32) ? 128'h00000000000000000000000080000000 :
				(tag == 33) ? 128'h00000000000000000000000100000000 :
				(tag == 34) ? 128'h00000000000000000000000200000000 :
				(tag == 35) ? 128'h00000000000000000000000400000000 :
				(tag == 36) ? 128'h00000000000000000000000800000000 :
				(tag == 37) ? 128'h00000000000000000000001000000000 :
				(tag == 38) ? 128'h00000000000000000000002000000000 :
				(tag == 39) ? 128'h00000000000000000000004000000000 :
				(tag == 40) ? 128'h00000000000000000000008000000000 :
				(tag == 41) ? 128'h00000000000000000000010000000000 :
				(tag == 42) ? 128'h00000000000000000000020000000000 :
				(tag == 43) ? 128'h00000000000000000000040000000000 :
				(tag == 44) ? 128'h00000000000000000000080000000000 :
				(tag == 45) ? 128'h00000000000000000000100000000000 :
				(tag == 46) ? 128'h00000000000000000000200000000000 :
				(tag == 47) ? 128'h00000000000000000000400000000000 :
				(tag == 48) ? 128'h00000000000000000000800000000000 :
				(tag == 49) ? 128'h00000000000000000001000000000000 :
				(tag == 50) ? 128'h00000000000000000002000000000000 :
				(tag == 51) ? 128'h00000000000000000004000000000000 :
				(tag == 52) ? 128'h00000000000000000008000000000000 :
				(tag == 53) ? 128'h00000000000000000010000000000000 :
				(tag == 54) ? 128'h00000000000000000020000000000000 :
				(tag == 55) ? 128'h00000000000000000040000000000000 :
				(tag == 56) ? 128'h00000000000000000080000000000000 :
				(tag == 57) ? 128'h00000000000000000100000000000000 :
				(tag == 58) ? 128'h00000000000000000200000000000000 :
				(tag == 59) ? 128'h00000000000000000400000000000000 :
				(tag == 60) ? 128'h00000000000000000800000000000000 :
				(tag == 61) ? 128'h00000000000000001000000000000000 :
				(tag == 62) ? 128'h00000000000000002000000000000000 :
				(tag == 63) ? 128'h00000000000000004000000000000000 :
				(tag == 64) ? 128'h00000000000000008000000000000000 :
				(tag == 65) ? 128'h00000000000000010000000000000000 :
				(tag == 66) ? 128'h00000000000000020000000000000000 :
				(tag == 67) ? 128'h00000000000000040000000000000000 :
				(tag == 68) ? 128'h00000000000000080000000000000000 :
				(tag == 69) ? 128'h00000000000000100000000000000000 :
				(tag == 70) ? 128'h00000000000000200000000000000000 :
				(tag == 71) ? 128'h00000000000000400000000000000000 :
				(tag == 72) ? 128'h00000000000000800000000000000000 :
				(tag == 73) ? 128'h00000000000001000000000000000000 :
				(tag == 74) ? 128'h00000000000002000000000000000000 :
				(tag == 75) ? 128'h00000000000004000000000000000000 :
				(tag == 76) ? 128'h00000000000008000000000000000000 :
				(tag == 77) ? 128'h00000000000010000000000000000000 :
				(tag == 78) ? 128'h00000000000020000000000000000000 :
				(tag == 79) ? 128'h00000000000040000000000000000000 :
				(tag == 80) ? 128'h00000000000080000000000000000000 :
				(tag == 81) ? 128'h00000000000100000000000000000000 :
				(tag == 82) ? 128'h00000000000200000000000000000000 :
				(tag == 83) ? 128'h00000000000400000000000000000000 :
				(tag == 84) ? 128'h00000000000800000000000000000000 :
				(tag == 85) ? 128'h00000000001000000000000000000000 :
				(tag == 86) ? 128'h00000000002000000000000000000000 :
				(tag == 87) ? 128'h00000000004000000000000000000000 :
				(tag == 88) ? 128'h00000000008000000000000000000000 :
				(tag == 89) ? 128'h00000000010000000000000000000000 :
				(tag == 90) ? 128'h00000000020000000000000000000000 :
				(tag == 91) ? 128'h00000000040000000000000000000000 :
				(tag == 92) ? 128'h00000000080000000000000000000000 :
				(tag == 93) ? 128'h00000000100000000000000000000000 :
				(tag == 94) ? 128'h00000000200000000000000000000000 :
				(tag == 95) ? 128'h00000000400000000000000000000000 :
				(tag == 96) ? 128'h00000000800000000000000000000000 :
				(tag == 97) ? 128'h00000001000000000000000000000000 :
				(tag == 98) ? 128'h00000002000000000000000000000000 :
				(tag == 99) ? 128'h00000004000000000000000000000000 :
				(tag == 100) ? 128'h00000008000000000000000000000000 :
				(tag == 101) ? 128'h00000010000000000000000000000000 :
				(tag == 102) ? 128'h00000020000000000000000000000000 :
				(tag == 103) ? 128'h00000040000000000000000000000000 :
				(tag == 104) ? 128'h00000080000000000000000000000000 :
				(tag == 105) ? 128'h00000100000000000000000000000000 :
				(tag == 106) ? 128'h00000200000000000000000000000000 :
				(tag == 107) ? 128'h00000400000000000000000000000000 :
				(tag == 108) ? 128'h00000800000000000000000000000000 :
				(tag == 109) ? 128'h00001000000000000000000000000000 :
				(tag == 110) ? 128'h00002000000000000000000000000000 :
				(tag == 111) ? 128'h00004000000000000000000000000000 :
				(tag == 112) ? 128'h00008000000000000000000000000000 :
				(tag == 113) ? 128'h00010000000000000000000000000000 :
				(tag == 114) ? 128'h00020000000000000000000000000000 :
				(tag == 115) ? 128'h00040000000000000000000000000000 :
				(tag == 116) ? 128'h00080000000000000000000000000000 :
				(tag == 117) ? 128'h00100000000000000000000000000000 :
				(tag == 118) ? 128'h00200000000000000000000000000000 :
				(tag == 119) ? 128'h00400000000000000000000000000000 :
				(tag == 120) ? 128'h00800000000000000000000000000000 :
				(tag == 121) ? 128'h01000000000000000000000000000000 :
				(tag == 122) ? 128'h02000000000000000000000000000000 :
				(tag == 123) ? 128'h04000000000000000000000000000000 :
				(tag == 124) ? 128'h08000000000000000000000000000000 :
				(tag == 125) ? 128'h10000000000000000000000000000000 :
				(tag == 126) ? 128'h20000000000000000000000000000000 :
				(tag == 127) ? 128'h40000000000000000000000000000000 :
				128'hxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;


endmodule