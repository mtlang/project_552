//Direct-mapped cache; 128 cache blocks
//Block # = (block address) % 128
//Above can be calculated by taking the low order 8 bits of address as block #
//The tag bits are the rest of the address not used for the index
//Word select bits are 3 least significant bits of the index
// i.e. index = address[7:0]
//      tag   = address[15:8]
//      word  = address[2:0]
module i_cache (clk, rst, Address, Data_In, Data_Out, Write_Enable, Miss);
input clk, rst, Write_Enable;
input [15:0] Address, Data_In;

output Miss;
output [15:0] Data_Out;

wire [2:0] word;
wire [7:0] tag_mda, tag, blk_index, word_en;
wire [15:0] cache_data;
wire [127:0] block_en;


//Decoder modules for one hot block enable and word enable
Decoder_7_128 dec_7_128(.tag(blk_index), .block(block_en));
decoder_3_8 dec_3_8(.A(word), .B(word_en));

//Meta data array (Valid + tag bits)
MetaDataArray MDA (.clk(clk), .rst(rst), .DataIn(tag), .Write(Write_Enable), .BlockEnable(block_en), .DataOut(tag_mda));

//Data array (cache lines)
DataArray DA (.clk(clk), .rst(rst), .DataIn(Data_In), .Write(Write_Enable), .BlockEnable(block_en), .WordEnable(word_en), .DataOut(cache_data));	

//first bit is valid bit in tag
assign tag = {1'b1,Address[14:8]};
assign blk_index = Address[7:0];
assign word = Address[2:0];

assign Miss = (~Write_Enable) ? (tag & tag_mda) : 1'b0;
assign Data_Out = (Write_Enable) ? 16'hxxxx : cache_data;

endmodule
